module main

fn main() {
	println('Mango - Compilador oficial v0.1.0-alpha')
}
